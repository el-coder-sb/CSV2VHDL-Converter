	--
	-- Measurement data of my_decoded_file.vhd starts here
	--
	wait for   0.0 ns;		spi_clk_stimu01_sl_s		<=	'1';
	wait for   0.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for 267.0 ns;		spi_mosi_stimu01_sl_s		<=	'1';
	wait for  24.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for  16.0 ns;		spi_mosi_stimu01_sl_s		<=	'1';
	wait for  38.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for  42.0 ns;		spi_mosi_stimu01_sl_s		<=	'1';
	wait for  38.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for  42.0 ns;		spi_mosi_stimu01_sl_s		<=	'1';
	wait for  24.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for 216.0 ns;		spi_mosi_stimu01_sl_s		<=	'1';
	wait for  24.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for  96.0 ns;		spi_mosi_stimu01_sl_s		<=	'1';
	wait for 163.0 ns;		spi_clk_stimu01_sl_s		<=	'0';
	wait for 440.0 ns;		spi_clk_stimu01_sl_s		<=	'1';
	wait for  20.0 ns;		spi_clk_stimu01_sl_s		<=	'0';
	wait for 825.0 ns;		spi_mosi_stimu01_sl_s		<=	'0';
	wait for  15.0 ns;		spi_clk_stimu01_sl_s		<=	'1';
